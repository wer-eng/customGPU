module DEMO_V01_TOP




endmodule
